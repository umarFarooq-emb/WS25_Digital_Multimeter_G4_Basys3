//  --------------------------------------------------------------------------
//                    Copyright Message
//  --------------------------------------------------------------------------
//
//  CONFIDENTIAL and PROPRIETARY
//  COPYRIGHT (c) XXXX 2019
//
//  All rights are reserved. Reproduction in whole or in part is
//  prohibited without the written consent of the copyright owner.
//
//
//  ----------------------------------------------------------------------------
//                    Design Information
//  ----------------------------------------------------------------------------
//
//  File             $URL: http://.../ste.sv $
//  Author
//  Date             $LastChangedDate: 2019-02-15 08:18:28 +0100 (Fri, 15 Feb 2019) $
//  Last changed by  $LastChangedBy: kstrohma $
//  Version          $Revision: 2472 $
//
// Description       Calculates the RMS value
//
//  ----------------------------------------------------------------------------
//                    Revision History (written manually)
//  ----------------------------------------------------------------------------
//
//  Date        Author     Change Description
//  ==========  =========  ========================================================
//  2019-01-09  strohmay   Initial verison       


// What is the limit in case I do a full calculation over the whole buffer after each sample
`default_nettype none
module ste_led_bar #(
  parameter int DATA_W                 =  4, 
  parameter logic[DATA_W-1:0] DATA_MAX =  1'hf,
  parameter int LED_NR                 =  8     // 
) (
  input   wire                clk             , // I; System clock 
  input   wire                rst_n           , // I; system cock reset (active low)  
  input   wire  [DATA_W-1:0]  din_i           , // I; Input data    
  input   wire                din_update_i    , // I; Input data update 
  input   wire                clr_i           , // I; Clear  data 
  output  logic [LED_NR-1:0]  led_o             // O; LEDs drive signal 
);
  
  
  // -------------------------------------------------------------------------
  // Definition 
  // -------------------------------------------------------------------------
  // make it big enough for multiplication later on
  logic [DATA_W+3:0] level;
    
  // -------------------------------------------------------------------------
  // Implementation
  // -------------------------------------------------------------------------

  // scale it to the be linear 
  //always_comb begin
  //  level = (din_i * LED_NR) / (DATA_MAX + 1);
  //end
    
 
  always_ff @(posedge clk) begin
    if (~rst_n || clr_i) begin
        led_o <= 0;
    end
    else if (din_update_i) begin
        // scale it to the be linear 
        level <= (din_i * LED_NR) / (DATA_MAX + 1);
        
        for (int i = 0; i < LED_NR; i++) begin
            led_o[i] <= (i <= level);
        end
    end
     
  end
  
endmodule

`default_nettype wire  